module rhythm_pcie (
);

endmodule